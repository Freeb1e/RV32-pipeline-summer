// Branch Target Buffer
// 用于建立PC值与分支指令及其分支地址之间的映射关系
module BTB(
        input wire clk,
        input wire rst,

        /* 时序逻辑， 更新buffer */
        input wire valid_in, // 是否有新的分支指令
        input wire [31:0] branch_PC, // 分支指令的PC值
        input wire [31:0] branch_target, // 分支指令的目标地址

        /* 组合逻辑 */
        input wire [31:0] PC_in, // 需要判断的PC值
        output wire is_branch_inst, // 是否为分支指令
        output wire [31:0] target_addr // 分支目标地址
    );

    // BTB参数定义
    parameter BTB_SIZE = 64;  // BTB表大小，必须是2的幂
    parameter INDEX_WIDTH = $clog2(BTB_SIZE);  // 索引位宽
    parameter TAG_WIDTH = 32 - INDEX_WIDTH - 2;  // 标签位宽 (PC - 索引位 - 字节偏移)

    // BTB表项定义
    reg [TAG_WIDTH-1:0] btb_tags [BTB_SIZE-1:0];  // 标签数组
    reg [31:0] btb_targets [BTB_SIZE-1:0];        // 目标地址数组
    reg btb_valid [BTB_SIZE-1:0];                 // 有效位数组

    // BTB索引计算 (使用PC的低位，忽略字节偏移)
    wire [INDEX_WIDTH-1:0] lookup_index = PC_in[INDEX_WIDTH+1:2];
    wire [TAG_WIDTH-1:0] lookup_tag = PC_in[31:INDEX_WIDTH+2];

    wire [INDEX_WIDTH-1:0] update_index = branch_PC[INDEX_WIDTH+1:2];
    wire [TAG_WIDTH-1:0] update_tag = branch_PC[31:INDEX_WIDTH+2];

    // 查找逻辑 - 判断当前PC是否命中BTB中的分支指令
    wire tag_match = (btb_tags[lookup_index] == lookup_tag);
    wire entry_valid = btb_valid[lookup_index];

    // 输出赋值
    assign is_branch_inst = tag_match && entry_valid;
    assign target_addr = (is_branch_inst) ? btb_targets[lookup_index] : 32'b0;

    // BTB更新逻辑
    integer i;
    always @(posedge clk) begin
        if (rst) begin
            // 复位时清空BTB表
            for (i = 0; i < BTB_SIZE; i = i + 1) begin
                btb_valid[i] <= 1'b0;
                btb_tags[i] <= {TAG_WIDTH{1'b0}};
                btb_targets[i] <= 32'b0;
            end
        end
        else if (valid_in) begin
            // 有新的分支指令时，更新BTB表
            btb_valid[update_index] <= 1'b1;
            btb_tags[update_index] <= update_tag;
            btb_targets[update_index] <= branch_target;
        end
    end

    // 未使用信号位注释
    // PC_in[1:0] 和 branch_PC[1:0] 未使用是正常的，因为是字节偏移
    /* verilator lint_off UNUSEDSIGNAL */

endmodule
